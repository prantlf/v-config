module config

import os { exists, getenv_opt, join_path_single, real_path }
import prantlf.debug { new_debug }

const d = new_debug('config')

const exts = [
	'.ini',
	'.properties',
	'.json',
	'.yml',
	'.yaml',
]!

pub fn find_config_file_any(start_dir string, name string, depth int, user bool) ?string {
	names := get_all_names(name)
	return find_config_file(start_dir, names, depth, user)
}

pub fn find_config_file(start_dir string, names []string, depth int, user bool) ?string {
	if config.d.is_enabled() {
		names_str := names.join('"", "')
		dstart_dir := config.d.rwd(start_dir)
		config.d.log_str('look for names "${names_str}" in "${dstart_dir}"')
	}

	mut dir := real_path(start_dir)
	for _ in -1 .. depth {
		file := find_file(dir, names)
		if file.len > 0 {
			return normalise_file(file)
		}
		dir = join_path_single(dir, '..')
	}

	if user {
		if home_dir := get_home_dir() {
			file := find_file(home_dir, names)
			if file.len > 0 {
				return normalise_file(file)
			}
		}
	}

	config.d.log_str('none of the names found')
	return none
}

pub fn find_user_config_file_any(name string) ?string {
	names := get_all_names(name)
	return find_user_config_file(names)
}

pub fn find_user_config_file(names []string) ?string {
	if home_dir := get_home_dir() {
		if config.d.is_enabled() {
			names_str := names.join('"", "')
			dhome_dir := config.d.rwd(home_dir)
			config.d.log_str('look for names "${names_str}" in "${dhome_dir}"')
		}

		file := find_file(home_dir, names)
		if file.len > 0 {
			return normalise_file(file)
		}

		config.d.log_str('none of the names found')
	}

	return none
}

fn normalise_file(path string) string {
	file := real_path(path)
	dfile := config.d.rwd(file)
	config.d.log('found "%s"', dfile)
	return file
}

fn find_file(dir string, names []string) string {
	for name in names {
		mut file := join_path_single(dir, name)
		mut ddir := config.d.rwd(dir)
		config.d.log('checking if "%s" exists in "%s"', name, ddir)
		if exists(file) {
			return file
		}
	}
	return ''
}

fn get_home_dir() ?string {
	var_name := $if windows {
		'USERPROFILE'
	} $else {
		'HOME'
	}
	return if home_dir := getenv_opt(var_name) {
		dhome_dir := config.d.rwd(home_dir)
		config.d.log('environment variable "%s" poins to "%s"', var_name, dhome_dir)
		home_dir
	} else {
		config.d.log('environment variable "%s" is empty', var_name)
		none
	}
}

fn get_all_names(name string) []string {
	mut names := []string{len: config.exts.len}
	for i in 0 .. config.exts.len {
		names[i] = '${name}${config.exts[i]}'
	}
	return names
}
